// Basic testbench for the SpeedPong game.

module speedPongTestbench();

endmodule